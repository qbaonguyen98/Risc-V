module ALU(alumux1_out, alumux2_out, aluop, aluout);
    input [31:0] alumux1_out, alumux2_out;
    input [3:0] aluop;

    output reg [31:0] aluout;

endmodule