module Reg();

endmodule